module secded_decoder (
  input  logic        CLK,
  input  logic [71:0] E_DATA,
  output logic [71:0] D_DATA,
  output logic        ERR,
  output logic        D_ERR,
  output logic        S_ERR
);

  logic [7:0]  SYNDROME;
  logic [71:0] MASK;
  logic        OR_SYND;
  logic        XOR_SYND;

  assign OR_SYND  = |SYNDROME;
  assign XOR_SYND = ^SYNDROME;

    // S1
    assign SYNDROME[0] = E_DATA[0] ^ E_DATA[1] ^ E_DATA[2] ^ E_DATA[3] ^ E_DATA[4] ^ E_DATA[5] ^ E_DATA[6] ^
	    E_DATA[7] ^ E_DATA[10] ^ E_DATA[13] ^ E_DATA[14] ^ E_DATA[17] ^ E_DATA[20] ^ E_DATA[23] ^
		  E_DATA[24] ^ E_DATA[27] ^ E_DATA[35] ^ E_DATA[43] ^ E_DATA[46] ^ E_DATA[47] ^ E_DATA[51] ^
		  E_DATA[52] ^ E_DATA[53] ^ E_DATA[56] ^ E_DATA[57] ^ E_DATA[58] ^ E_DATA[64];
    
    // S2
    assign SYNDROME[1] = E_DATA[0] ^ E_DATA[1] ^ E_DATA[2] ^ E_DATA[8] ^ E_DATA[9] ^ E_DATA[10] ^ E_DATA[11] ^
	    E_DATA[12] ^ E_DATA[13] ^ E_DATA[14] ^ E_DATA[15] ^ E_DATA[18] ^ E_DATA[21] ^ E_DATA[22] ^
		  E_DATA[25] ^ E_DATA[28] ^ E_DATA[31] ^ E_DATA[32] ^ E_DATA[35] ^ E_DATA[43] ^ E_DATA[51] ^
		  E_DATA[54] ^ E_DATA[55] ^ E_DATA[59] ^ E_DATA[60] ^ E_DATA[61] ^ E_DATA[65];

    // S3
    assign SYNDROME[2] = E_DATA[3] ^ E_DATA[4] ^ E_DATA[5] ^ E_DATA[8] ^ E_DATA[9] ^ E_DATA[10] ^ E_DATA[16] ^
	    E_DATA[17] ^ E_DATA[18] ^ E_DATA[19] ^ E_DATA[20] ^ E_DATA[21] ^ E_DATA[22] ^ E_DATA[23] ^
		  E_DATA[26] ^ E_DATA[29] ^ E_DATA[30] ^ E_DATA[33] ^ E_DATA[36] ^ E_DATA[39] ^ E_DATA[40] ^
		  E_DATA[43] ^ E_DATA[51] ^ E_DATA[59] ^ E_DATA[62] ^ E_DATA[63] ^ E_DATA[66];

    // S4
    assign SYNDROME[3] = E_DATA[3] ^ E_DATA[6] ^ E_DATA[7] ^ E_DATA[11] ^ E_DATA[12] ^ E_DATA[13] ^ E_DATA[16] ^ 
		  E_DATA[17] ^ E_DATA[18] ^ E_DATA[24] ^ E_DATA[25] ^ E_DATA[26] ^ E_DATA[27] ^ E_DATA[28] ^ 
		  E_DATA[29] ^ E_DATA[30] ^ E_DATA[31] ^ E_DATA[34] ^ E_DATA[37] ^ E_DATA[38] ^ E_DATA[41] ^ 
		  E_DATA[44] ^ E_DATA[47] ^ E_DATA[48] ^ E_DATA[51] ^ E_DATA[59] ^ E_DATA[67];

    // S5
    assign SYNDROME[4] = E_DATA[3] ^ E_DATA[11] ^ E_DATA[14] ^ E_DATA[15] ^ E_DATA[19] ^ E_DATA[20] ^ E_DATA[21] ^
	    E_DATA[24] ^ E_DATA[25] ^ E_DATA[26] ^ E_DATA[32] ^ E_DATA[33] ^ E_DATA[34] ^ E_DATA[35] ^
		  E_DATA[36] ^ E_DATA[37] ^ E_DATA[38] ^ E_DATA[39] ^ E_DATA[42] ^ E_DATA[45] ^ E_DATA[46] ^
		  E_DATA[49] ^ E_DATA[52] ^ E_DATA[55] ^ E_DATA[56] ^ E_DATA[59] ^ E_DATA[68];

    // S6
    assign SYNDROME[5] = E_DATA[0] ^ E_DATA[3] ^ E_DATA[11] ^ E_DATA[19] ^ E_DATA[22] ^ E_DATA[23] ^ E_DATA[27] ^
	    E_DATA[28] ^ E_DATA[29] ^ E_DATA[32] ^ E_DATA[33] ^ E_DATA[34] ^ E_DATA[40] ^ E_DATA[41] ^
		  E_DATA[42] ^ E_DATA[43] ^ E_DATA[44] ^ E_DATA[45] ^ E_DATA[46] ^ E_DATA[47] ^ E_DATA[50] ^
		  E_DATA[53] ^ E_DATA[54] ^ E_DATA[57] ^ E_DATA[60] ^ E_DATA[63] ^ E_DATA[69];

    // S7
    assign SYNDROME[6] = E_DATA[1] ^ E_DATA[4] ^ E_DATA[7] ^ E_DATA[8] ^ E_DATA[11] ^ E_DATA[19] ^ E_DATA[27] ^
	    E_DATA[30] ^ E_DATA[31] ^ E_DATA[35] ^ E_DATA[36] ^ E_DATA[37] ^ E_DATA[40] ^ E_DATA[41] ^
		  E_DATA[42] ^ E_DATA[48] ^ E_DATA[49] ^ E_DATA[50] ^ E_DATA[51] ^ E_DATA[52] ^ E_DATA[53] ^
		  E_DATA[54] ^ E_DATA[55] ^ E_DATA[58] ^ E_DATA[61] ^ E_DATA[62] ^ E_DATA[70];

    // S8
    assign SYNDROME[7] = E_DATA[2] ^ E_DATA[5] ^ E_DATA[6] ^ E_DATA[9] ^ E_DATA[12] ^ E_DATA[15] ^ E_DATA[16] ^
	    E_DATA[19] ^ E_DATA[27] ^ E_DATA[35] ^ E_DATA[38] ^ E_DATA[39] ^ E_DATA[43] ^ E_DATA[44] ^
		  E_DATA[45] ^ E_DATA[48] ^ E_DATA[49] ^ E_DATA[50] ^ E_DATA[56] ^ E_DATA[57] ^ E_DATA[58] ^
		  E_DATA[59] ^ E_DATA[60] ^ E_DATA[61] ^ E_DATA[62] ^ E_DATA[63] ^ E_DATA[71];

  always @(posedge CLK) begin
    ERR      <= OR_SYND;
    D_ERR    <= OR_SYND & !XOR_SYND;
    S_ERR    <= OR_SYND & XOR_SYND;
    D_DATA   <= MASK ^ E_DATA;
    
  end

  always @(*) begin
    case (SYNDROME) 
      8'b00100011: MASK = 72'h00_0000_0000_0000_0001; // E_DATA[0]
      8'b01000011: MASK = 72'h00_0000_0000_0000_0002; // E_DATA[1]
      8'b10000011: MASK = 72'h00_0000_0000_0000_0004; // E_DATA[2]
      8'b00111101: MASK = 72'h00_0000_0000_0000_0008; // E_DATA[3]
      8'b01000101: MASK = 72'h00_0000_0000_0000_0010; // E_DATA[4]
      8'b10000101: MASK = 72'h00_0000_0000_0000_0020; // E_DATA[5]
      8'b10001001: MASK = 72'h00_0000_0000_0000_0040; // E_DATA[6]
      8'b01001001: MASK = 72'h00_0000_0000_0000_0080; // E_DATA[7]
      8'b01000110: MASK = 72'h00_0000_0000_0000_0100; // E_DATA[8]
      8'b10000110: MASK = 72'h00_0000_0000_0000_0200; // E_DATA[9]
      8'b00000111: MASK = 72'h00_0000_0000_0000_0400; // E_DATA[10]
      8'b01111010: MASK = 72'h00_0000_0000_0000_0800; // E_DATA[11]
      8'b10001010: MASK = 72'h00_0000_0000_0000_1000; // E_DATA[12]
      8'b00001011: MASK = 72'h00_0000_0000_0000_2000; // E_DATA[13]
      8'b00010011: MASK = 72'h00_0000_0000_0000_4000; // E_DATA[14]
      8'b10010010: MASK = 72'h00_0000_0000_0000_8000; // E_DATA[15]
      8'b10001100: MASK = 72'h00_0000_0000_0001_0000; // E_DATA[16]
      8'b00001101: MASK = 72'h00_0000_0000_0002_0000; // E_DATA[17]
      8'b00001110: MASK = 72'h00_0000_0000_0004_0000; // E_DATA[18]
      8'b11110100: MASK = 72'h00_0000_0000_0008_0000; // E_DATA[19]
      8'b00010101: MASK = 72'h00_0000_0000_0010_0000; // E_DATA[20]
      8'b00010110: MASK = 72'h00_0000_0000_0020_0000; // E_DATA[21]
      8'b00100110: MASK = 72'h00_0000_0000_0040_0000; // E_DATA[22]
      8'b00100101: MASK = 72'h00_0000_0000_0080_0000; // E_DATA[23]
      8'b00011001: MASK = 72'h00_0000_0000_0100_0000; // E_DATA[24]
      8'b00011010: MASK = 72'h00_0000_0000_0200_0000; // E_DATA[25]
      8'b00011100: MASK = 72'h00_0000_0000_0400_0000; // E_DATA[26]
      8'b11101001: MASK = 72'h00_0000_0000_0800_0000; // E_DATA[27]
      8'b00101010: MASK = 72'h00_0000_0000_1000_0000; // E_DATA[28]
      8'b00101100: MASK = 72'h00_0000_0000_2000_0000; // E_DATA[29]
      8'b01001100: MASK = 72'h00_0000_0000_4000_0000; // E_DATA[30]
      8'b01001010: MASK = 72'h00_0000_0000_8000_0000; // E_DATA[31]
      8'b00110010: MASK = 72'h00_0000_0001_0000_0000; // E_DATA[32]
      8'b00110100: MASK = 72'h00_0000_0002_0000_0000; // E_DATA[33]
      8'b00111000: MASK = 72'h00_0000_0004_0000_0000; // E_DATA[34]
      8'b11010011: MASK = 72'h00_0000_0008_0000_0000; // E_DATA[35]
      8'b01010100: MASK = 72'h00_0000_0010_0000_0000; // E_DATA[36]
      8'b01011000: MASK = 72'h00_0000_0020_0000_0000; // E_DATA[37]
      8'b10011000: MASK = 72'h00_0000_0040_0000_0000; // E_DATA[38]
      8'b10010100: MASK = 72'h00_0000_0080_0000_0000; // E_DATA[39]
      8'b01100100: MASK = 72'h00_0000_0100_0000_0000; // E_DATA[40]
      8'b01101000: MASK = 72'h00_0000_0200_0000_0000; // E_DATA[41]
      8'b01110000: MASK = 72'h00_0000_0400_0000_0000; // E_DATA[42]
      8'b10100111: MASK = 72'h00_0000_0800_0000_0000; // E_DATA[43]
      8'b10101000: MASK = 72'h00_0000_1000_0000_0000; // E_DATA[44]
      8'b10110000: MASK = 72'h00_0000_2000_0000_0000; // E_DATA[45]
      8'b00110001: MASK = 72'h00_0000_4000_0000_0000; // E_DATA[46]
      8'b00101001: MASK = 72'h00_0000_8000_0000_0000; // E_DATA[47]
      8'b11001000: MASK = 72'h00_0001_0000_0000_0000; // E_DATA[48]
      8'b11010000: MASK = 72'h00_0002_0000_0000_0000; // E_DATA[49]
      8'b11100000: MASK = 72'h00_0004_0000_0000_0000; // E_DATA[50]
      8'b01001111: MASK = 72'h00_0008_0000_0000_0000; // E_DATA[51]
      8'b01010001: MASK = 72'h00_0010_0000_0000_0000; // E_DATA[52]
      8'b01100001: MASK = 72'h00_0020_0000_0000_0000; // E_DATA[53]
      8'b01100010: MASK = 72'h00_0040_0000_0000_0000; // E_DATA[54]
      8'b01010010: MASK = 72'h00_0080_0000_0000_0000; // E_DATA[55]
      8'b10010001: MASK = 72'h00_0100_0000_0000_0000; // E_DATA[56]
      8'b10100001: MASK = 72'h00_0200_0000_0000_0000; // E_DATA[57]
      8'b11000001: MASK = 72'h00_0400_0000_0000_0000; // E_DATA[58]
      8'b10011110: MASK = 72'h00_0800_0000_0000_0000; // E_DATA[59]
      8'b10100010: MASK = 72'h00_1000_0000_0000_0000; // E_DATA[60]
      8'b11000010: MASK = 72'h00_2000_0000_0000_0000; // E_DATA[61]
      8'b11000100: MASK = 72'h00_4000_0000_0000_0000; // E_DATA[62]
      8'b10100100: MASK = 72'h00_8000_0000_0000_0000; // E_DATA[63]
      8'b00000001: MASK = 72'h01_0000_0000_0000_0000; // E_DATA[64]
      8'b00000010: MASK = 72'h02_0000_0000_0000_0000; // E_DATA[65]
      8'b00000100: MASK = 72'h04_0000_0000_0000_0000; // E_DATA[66]
      8'b00001000: MASK = 72'h08_0000_0000_0000_0000; // E_DATA[67]
      8'b00010000: MASK = 72'h10_0000_0000_0000_0000; // E_DATA[68]
      8'b00100000: MASK = 72'h20_0000_0000_0000_0000; // E_DATA[69]
      8'b01000000: MASK = 72'h40_0000_0000_0000_0000; // E_DATA[70]
      8'b10000000: MASK = 72'h80_0000_0000_0000_0000; // E_DATA[71]
      default:     MASK = 72'h00_0000_0000_0000_0000; // no error
    endcase
   end
endmodule
