module secded_decoder (
  input  logic        CLK,
  input  logic [71:0] E_DATA,
  output logic [71:0] D_DATA,
  output logic        ERR,
  output logic        D_ERR,
  output logic        S_ERR
);

  logic [71:0] BUFFER;
  logic [7:0]  SYNDROME;
  logic [71:0] MASK;
  logic        OR_SYND;
  logic        XOR_SYND;

  assign OR_SYND  = |SYNDROME;
  assign XOR_SYND = ^SYNDROME;
  assign ERR      = OR_SYND;
  assign D_ERR    = OR_SYND & !XOR_SYND;
  assign S_ERR    = OR_SYND & XOR_SYND;
  assign D_DATA   = MASK ^ BUFFER;
    
  // S1
  assign SYNDROME[0] = BUFFER[0] ^ BUFFER[1] ^ BUFFER[2] ^ BUFFER[3] ^ BUFFER[4] ^ BUFFER[5] ^ BUFFER[6] ^
	  BUFFER[7] ^ BUFFER[10] ^ BUFFER[13] ^ BUFFER[14] ^ BUFFER[17] ^ BUFFER[20] ^ BUFFER[23] ^
		BUFFER[24] ^ BUFFER[27] ^ BUFFER[35] ^ BUFFER[43] ^ BUFFER[46] ^ BUFFER[47] ^ BUFFER[51] ^
		BUFFER[52] ^ BUFFER[53] ^ BUFFER[56] ^ BUFFER[57] ^ BUFFER[58] ^ BUFFER[64];
    
  // S2
  assign SYNDROME[1] = BUFFER[0] ^ BUFFER[1] ^ BUFFER[2] ^ BUFFER[8] ^ BUFFER[9] ^ BUFFER[10] ^ BUFFER[11] ^
	  BUFFER[12] ^ BUFFER[13] ^ BUFFER[14] ^ BUFFER[15] ^ BUFFER[18] ^ BUFFER[21] ^ BUFFER[22] ^
		BUFFER[25] ^ BUFFER[28] ^ BUFFER[31] ^ BUFFER[32] ^ BUFFER[35] ^ BUFFER[43] ^ BUFFER[51] ^
		BUFFER[54] ^ BUFFER[55] ^ BUFFER[59] ^ BUFFER[60] ^ BUFFER[61] ^ BUFFER[65];

  // S3
  assign SYNDROME[2] = BUFFER[3] ^ BUFFER[4] ^ BUFFER[5] ^ BUFFER[8] ^ BUFFER[9] ^ BUFFER[10] ^ BUFFER[16] ^
    BUFFER[17] ^ BUFFER[18] ^ BUFFER[19] ^ BUFFER[20] ^ BUFFER[21] ^ BUFFER[22] ^ BUFFER[23] ^
    BUFFER[26] ^ BUFFER[29] ^ BUFFER[30] ^ BUFFER[33] ^ BUFFER[36] ^ BUFFER[39] ^ BUFFER[40] ^
    BUFFER[43] ^ BUFFER[51] ^ BUFFER[59] ^ BUFFER[62] ^ BUFFER[63] ^ BUFFER[66];

    // S4
  assign SYNDROME[3] = BUFFER[3] ^ BUFFER[6] ^ BUFFER[7] ^ BUFFER[11] ^ BUFFER[12] ^ BUFFER[13] ^ BUFFER[16] ^ 
		BUFFER[17] ^ BUFFER[18] ^ BUFFER[24] ^ BUFFER[25] ^ BUFFER[26] ^ BUFFER[27] ^ BUFFER[28] ^ 
		BUFFER[29] ^ BUFFER[30] ^ BUFFER[31] ^ BUFFER[34] ^ BUFFER[37] ^ BUFFER[38] ^ BUFFER[41] ^ 
		BUFFER[44] ^ BUFFER[47] ^ BUFFER[48] ^ BUFFER[51] ^ BUFFER[59] ^ BUFFER[67];

  // S5
  assign SYNDROME[4] = BUFFER[3] ^ BUFFER[11] ^ BUFFER[14] ^ BUFFER[15] ^ BUFFER[19] ^ BUFFER[20] ^ BUFFER[21] ^
    BUFFER[24] ^ BUFFER[25] ^ BUFFER[26] ^ BUFFER[32] ^ BUFFER[33] ^ BUFFER[34] ^ BUFFER[35] ^
	  BUFFER[36] ^ BUFFER[37] ^ BUFFER[38] ^ BUFFER[39] ^ BUFFER[42] ^ BUFFER[45] ^ BUFFER[46] ^
	  BUFFER[49] ^ BUFFER[52] ^ BUFFER[55] ^ BUFFER[56] ^ BUFFER[59] ^ BUFFER[68];

  // S6
  assign SYNDROME[5] = BUFFER[0] ^ BUFFER[3] ^ BUFFER[11] ^ BUFFER[19] ^ BUFFER[22] ^ BUFFER[23] ^ BUFFER[27] ^
    BUFFER[28] ^ BUFFER[29] ^ BUFFER[32] ^ BUFFER[33] ^ BUFFER[34] ^ BUFFER[40] ^ BUFFER[41] ^
	  BUFFER[42] ^ BUFFER[43] ^ BUFFER[44] ^ BUFFER[45] ^ BUFFER[46] ^ BUFFER[47] ^ BUFFER[50] ^
	  BUFFER[53] ^ BUFFER[54] ^ BUFFER[57] ^ BUFFER[60] ^ BUFFER[63] ^ BUFFER[69];

  // S7
  assign SYNDROME[6] = BUFFER[1] ^ BUFFER[4] ^ BUFFER[7] ^ BUFFER[8] ^ BUFFER[11] ^ BUFFER[19] ^ BUFFER[27] ^
    BUFFER[30] ^ BUFFER[31] ^ BUFFER[35] ^ BUFFER[36] ^ BUFFER[37] ^ BUFFER[40] ^ BUFFER[41] ^
	  BUFFER[42] ^ BUFFER[48] ^ BUFFER[49] ^ BUFFER[50] ^ BUFFER[51] ^ BUFFER[52] ^ BUFFER[53] ^
	  BUFFER[54] ^ BUFFER[55] ^ BUFFER[58] ^ BUFFER[61] ^ BUFFER[62] ^ BUFFER[70];

  // S8
  assign SYNDROME[7] = BUFFER[2] ^ BUFFER[5] ^ BUFFER[6] ^ BUFFER[9] ^ BUFFER[12] ^ BUFFER[15] ^ BUFFER[16] ^
    BUFFER[19] ^ BUFFER[27] ^ BUFFER[35] ^ BUFFER[38] ^ BUFFER[39] ^ BUFFER[43] ^ BUFFER[44] ^
	  BUFFER[45] ^ BUFFER[48] ^ BUFFER[49] ^ BUFFER[50] ^ BUFFER[56] ^ BUFFER[57] ^ BUFFER[58] ^
	  BUFFER[59] ^ BUFFER[60] ^ BUFFER[61] ^ BUFFER[62] ^ BUFFER[63] ^ BUFFER[71];

  always @(posedge CLK) begin
    BUFFER <= E_DATA;
  end

  always @(*) begin
    case (SYNDROME) 
      8'b00100011: MASK = 72'h00_0000_0000_0000_0001; // BUFFER[0]
      8'b01000011: MASK = 72'h00_0000_0000_0000_0002; // BUFFER[1]
      8'b10000011: MASK = 72'h00_0000_0000_0000_0004; // BUFFER[2]
      8'b00111101: MASK = 72'h00_0000_0000_0000_0008; // BUFFER[3]
      8'b01000101: MASK = 72'h00_0000_0000_0000_0010; // BUFFER[4]
      8'b10000101: MASK = 72'h00_0000_0000_0000_0020; // BUFFER[5]
      8'b10001001: MASK = 72'h00_0000_0000_0000_0040; // BUFFER[6]
      8'b01001001: MASK = 72'h00_0000_0000_0000_0080; // BUFFER[7]
      8'b01000110: MASK = 72'h00_0000_0000_0000_0100; // BUFFER[8]
      8'b10000110: MASK = 72'h00_0000_0000_0000_0200; // BUFFER[9]
      8'b00000111: MASK = 72'h00_0000_0000_0000_0400; // BUFFER[10]
      8'b01111010: MASK = 72'h00_0000_0000_0000_0800; // BUFFER[11]
      8'b10001010: MASK = 72'h00_0000_0000_0000_1000; // BUFFER[12]
      8'b00001011: MASK = 72'h00_0000_0000_0000_2000; // BUFFER[13]
      8'b00010011: MASK = 72'h00_0000_0000_0000_4000; // BUFFER[14]
      8'b10010010: MASK = 72'h00_0000_0000_0000_8000; // BUFFER[15]
      8'b10001100: MASK = 72'h00_0000_0000_0001_0000; // BUFFER[16]
      8'b00001101: MASK = 72'h00_0000_0000_0002_0000; // BUFFER[17]
      8'b00001110: MASK = 72'h00_0000_0000_0004_0000; // BUFFER[18]
      8'b11110100: MASK = 72'h00_0000_0000_0008_0000; // BUFFER[19]
      8'b00010101: MASK = 72'h00_0000_0000_0010_0000; // BUFFER[20]
      8'b00010110: MASK = 72'h00_0000_0000_0020_0000; // BUFFER[21]
      8'b00100110: MASK = 72'h00_0000_0000_0040_0000; // BUFFER[22]
      8'b00100101: MASK = 72'h00_0000_0000_0080_0000; // BUFFER[23]
      8'b00011001: MASK = 72'h00_0000_0000_0100_0000; // BUFFER[24]
      8'b00011010: MASK = 72'h00_0000_0000_0200_0000; // BUFFER[25]
      8'b00011100: MASK = 72'h00_0000_0000_0400_0000; // BUFFER[26]
      8'b11101001: MASK = 72'h00_0000_0000_0800_0000; // BUFFER[27]
      8'b00101010: MASK = 72'h00_0000_0000_1000_0000; // BUFFER[28]
      8'b00101100: MASK = 72'h00_0000_0000_2000_0000; // BUFFER[29]
      8'b01001100: MASK = 72'h00_0000_0000_4000_0000; // BUFFER[30]
      8'b01001010: MASK = 72'h00_0000_0000_8000_0000; // BUFFER[31]
      8'b00110010: MASK = 72'h00_0000_0001_0000_0000; // BUFFER[32]
      8'b00110100: MASK = 72'h00_0000_0002_0000_0000; // BUFFER[33]
      8'b00111000: MASK = 72'h00_0000_0004_0000_0000; // BUFFER[34]
      8'b11010011: MASK = 72'h00_0000_0008_0000_0000; // BUFFER[35]
      8'b01010100: MASK = 72'h00_0000_0010_0000_0000; // BUFFER[36]
      8'b01011000: MASK = 72'h00_0000_0020_0000_0000; // BUFFER[37]
      8'b10011000: MASK = 72'h00_0000_0040_0000_0000; // BUFFER[38]
      8'b10010100: MASK = 72'h00_0000_0080_0000_0000; // BUFFER[39]
      8'b01100100: MASK = 72'h00_0000_0100_0000_0000; // BUFFER[40]
      8'b01101000: MASK = 72'h00_0000_0200_0000_0000; // BUFFER[41]
      8'b01110000: MASK = 72'h00_0000_0400_0000_0000; // BUFFER[42]
      8'b10100111: MASK = 72'h00_0000_0800_0000_0000; // BUFFER[43]
      8'b10101000: MASK = 72'h00_0000_1000_0000_0000; // BUFFER[44]
      8'b10110000: MASK = 72'h00_0000_2000_0000_0000; // BUFFER[45]
      8'b00110001: MASK = 72'h00_0000_4000_0000_0000; // BUFFER[46]
      8'b00101001: MASK = 72'h00_0000_8000_0000_0000; // BUFFER[47]
      8'b11001000: MASK = 72'h00_0001_0000_0000_0000; // BUFFER[48]
      8'b11010000: MASK = 72'h00_0002_0000_0000_0000; // BUFFER[49]
      8'b11100000: MASK = 72'h00_0004_0000_0000_0000; // BUFFER[50]
      8'b01001111: MASK = 72'h00_0008_0000_0000_0000; // BUFFER[51]
      8'b01010001: MASK = 72'h00_0010_0000_0000_0000; // BUFFER[52]
      8'b01100001: MASK = 72'h00_0020_0000_0000_0000; // BUFFER[53]
      8'b01100010: MASK = 72'h00_0040_0000_0000_0000; // BUFFER[54]
      8'b01010010: MASK = 72'h00_0080_0000_0000_0000; // BUFFER[55]
      8'b10010001: MASK = 72'h00_0100_0000_0000_0000; // BUFFER[56]
      8'b10100001: MASK = 72'h00_0200_0000_0000_0000; // BUFFER[57]
      8'b11000001: MASK = 72'h00_0400_0000_0000_0000; // BUFFER[58]
      8'b10011110: MASK = 72'h00_0800_0000_0000_0000; // BUFFER[59]
      8'b10100010: MASK = 72'h00_1000_0000_0000_0000; // BUFFER[60]
      8'b11000010: MASK = 72'h00_2000_0000_0000_0000; // BUFFER[61]
      8'b11000100: MASK = 72'h00_4000_0000_0000_0000; // BUFFER[62]
      8'b10100100: MASK = 72'h00_8000_0000_0000_0000; // BUFFER[63]
      8'b00000001: MASK = 72'h01_0000_0000_0000_0000; // BUFFER[64]
      8'b00000010: MASK = 72'h02_0000_0000_0000_0000; // BUFFER[65]
      8'b00000100: MASK = 72'h04_0000_0000_0000_0000; // BUFFER[66]
      8'b00001000: MASK = 72'h08_0000_0000_0000_0000; // BUFFER[67]
      8'b00010000: MASK = 72'h10_0000_0000_0000_0000; // BUFFER[68]
      8'b00100000: MASK = 72'h20_0000_0000_0000_0000; // BUFFER[69]
      8'b01000000: MASK = 72'h40_0000_0000_0000_0000; // BUFFER[70]
      8'b10000000: MASK = 72'h80_0000_0000_0000_0000; // BUFFER[71]
      default:     MASK = 72'h00_0000_0000_0000_0000; // no error
    endcase
   end
endmodule
